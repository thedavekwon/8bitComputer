module mux2to1(din1, din2, dout);
   
   input din1, din2;
   output dout;

endmodule

module mux4to1(din1, din2, din3, din4,  dout);
   
   input din1, din2, din3, din4;
   output dout;

endmodule
