module shiftregs(din, dout, select);
   
   input [7:0] din;
   input       select;
   output [7:0] dout;
   
  
endmodule
