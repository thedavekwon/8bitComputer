module pc(din, dout);
   
   input din;
   output dout;
   
  
endmodule
