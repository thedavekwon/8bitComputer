module alu (instruction, acc, regIn, regOut);
   
	input [7:0] instruction, acc, regIn;
	output [7:0] regOut;
   
endmodule 
