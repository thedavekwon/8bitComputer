module controlunit(instruction, dout1, dout2, dout3);
   
   input instruction;
   output [7:0] dout1. dout2, dout3;
   
  
endmodule
